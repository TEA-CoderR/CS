module ptw {
	input clk;
	input rst;

	//TLB Interface
	input 
};